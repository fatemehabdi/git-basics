
Git Basics
-------------
I am learning the basics of git and github so 