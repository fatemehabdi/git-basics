---title new code 
---- new project accelleration
entity 

end; 

Git Basics
-------------

 
if a> basics
 c <= a+b ; 
then 

while 1 = abs
 end 
if  a> 1 then 
end
 
 -- chenges in github site 

