
Git Basics
-------------
I am learning the basics of git and github so 

if a> basics
else c = 2
then 
