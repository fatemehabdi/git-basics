---title new code 
---- new project accelleration
entity 
port(a in )
end; 

Git Basics
-------------
I am learning the basics of git and github so 

if a> basics
else c = 2
then 

while 1 = abs

if e 
else 
end

