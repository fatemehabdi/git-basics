---title new code 
---- new project accelleration
entity 
port(a in )
end; 

Git Basics
-------------
-- new changes in code 
 
if a> basics

then 

while 1 = abs
 end 
if  a> 1 then 
else 
end

